library verilog;
use verilog.vl_types.all;
entity UART_RX_tb is
end UART_RX_tb;
